`timescale 1ns / 1ps



module pingpong_test;
reg CLK,RST_N,FILP,HOLD;
wire [4:0] OUT;
wire DIR,MIN,MAX;

pingpong pp1(CLK,RST_N,OUT,MAX,MIN,HOLD,FILP,DIR);

initial begin
$fsdbDumpfile("Majority.fsdb");
$fsdbDumpvars;
end 

initial begin //initialization
//--------------------------------------------------------------------------------------------------------------------------
#0 CLK <= 1'b0; RST_N <= 1'b0; HOLD <= 1'b0; FILP <= 1'b0;
//Start running
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; 
//Single Variable (Fit with clk)
//--------------------------------------------------------------------------------------------------------------------------
#350 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b0; //Reset triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Rest triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b0; //Hold triggered on  
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b1; //Filp triggered on (one clock)
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b1; // Filp triggered on (multi clock) 
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b0; //Filp triggered off
//Double Variables (Fit with clk)
//-------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //initialization
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b0; HOLD = 1'b1; FILP = 1'b0; //Reset & Hold triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Reset & Hold triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b1; //Reset & Filp triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Reset & Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b1; //Hold & Filp triggered on(one clk)
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold & Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b1; //Hold & Filp triggered on(multi clk)
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold & Filp triggered off
//Single Variable(Asynthesize)
//--------------------------------------------------------------------------------------------------------------------------
#51 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b0; //Reset triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Rest triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b0; //Hold triggered on  
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold triggered off
//--------------------------------------------------------------------------------------------------------------------------
#18 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b1; //Filp triggered on (one clock)
//--------------------------------------------------------------------------------------------------------------------------
#32 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b1; // Filp triggered on (multi clock) 
//--------------------------------------------------------------------------------------------------------------------------
#59 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b0; //Filp triggered off
//Double Variables (Asynthesize)
//--------------------------------------------------------------------------------------------------------------------------
#51 RST_N = 1'b0; HOLD = 1'b1; FILP = 1'b0; //Reset & Hold triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Reset & Hold triggered off
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b0; HOLD = 1'b0; FILP = 1'b1; //Reset & Filp triggered on
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Reset & Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#18 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b1; //Hold & Filp triggered on(one clk)
//--------------------------------------------------------------------------------------------------------------------------
#32 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold & Filp triggered off
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b1; HOLD = 1'b1; FILP = 1'b1; //Hold & Filp triggered on(multi clk)
//--------------------------------------------------------------------------------------------------------------------------
#59 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; //Hold & Filp triggered off
//All variable
//--------------------------------------------------------------------------------------------------------------------------
#50 RST_N = 1'b0; HOLD = 1'b1; FILP = 1'b1; //Reset&Hold & Filp triggered on
//initialation
//--------------------------------------------------------------------------------------------------------------------------
#10 RST_N = 1'b1; HOLD = 1'b0; FILP = 1'b0; 
//--------------------------------------------------------------------------------------------------------------------------
end
//clk setting
always #5 CLK <= ~CLK;
//Termination condition
initial 
begin
#5000 $finish;
end
endmodule


